** Profile: "SCHEMATIC1-series"  [ E:\orcad\Regulator_circuit\Series_voltage_regulator_circuit-PSpiceFiles\SCHEMATIC1\series.sim ] 

** Creating circuit file "series.cir" 
** WARNING: THIS AUTOMATICALLY GENERATED FILE MAY BE OVERWRITTEN BY SUBSEQUENT SIMULATIONS

*Libraries: 
* Profile Libraries :
* Local Libraries :
* From [PSPICE NETLIST] section of C:\SPB_Data\cdssetup\OrCAD_PSpice\17.2.0\PSpice.ini file:
.lib "nomd.lib" 

*Analysis directives: 
.TRAN  0 200ms 0 
.STEP PARAM amp LIST 100,300,380,500,50000 
.OPTIONS ADVCONV
.PROBE64 V(alias(*)) I(alias(*)) W(alias(*)) D(alias(*)) NOISE(alias(*)) 
.INC "..\SCHEMATIC1.net" 


.END
